
// Code your design here
module ex;
  int i;
  initial begin
    while(i<=10)begin
      $display("value of i = %0d",i);
      i++;
    end
  end
endmodule


# value of i = 0
# value of i = 1
# value of i = 2
# value of i = 3
# value of i = 4
# value of i = 5
# value of i = 6
# value of i = 7
# value of i = 8
# value of i = 9
# value of i = 10
