module exam;
  int i;
  initial begin
    for(int i=0; i<=10; i++)
      $display("The Value Of i =%0d",i);
    
  end
endmodule


# The Value Of i =0
# The Value Of i =1
# The Value Of i =2
# The Value Of i =3
# The Value Of i =4
# The Value Of i =5
# The Value Of i =6
# The Value Of i =7
# The Value Of i =8
# The Value Of i =9
# The Value Of i =10
