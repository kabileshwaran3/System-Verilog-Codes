module mixed_array;
  reg [3:0][2:0]data[2:0][4:0];
  initial begin
    foreach(data[i,j,k,l])begin
      data[i][j][k][l]=$random;
      $display("Mixed Array data[%0d][%0d][%0d][%0d]=%d",i,j,k,l,data[i][j][k][l]);
    end
  end
    
endmodule                 
                    
                

output
# Mixed Array data[2][4][3][2]=0
# Mixed Array data[2][4][3][1]=1
# Mixed Array data[2][4][3][0]=1
# Mixed Array data[2][4][2][2]=1
# Mixed Array data[2][4][2][1]=1
# Mixed Array data[2][4][2][0]=1
# Mixed Array data[2][4][1][2]=1
# Mixed Array data[2][4][1][1]=0
# Mixed Array data[2][4][1][0]=1
# Mixed Array data[2][4][0][2]=1
# Mixed Array data[2][4][0][1]=0
# Mixed Array data[2][4][0][0]=1
# Mixed Array data[2][3][3][2]=1
# Mixed Array data[2][3][3][1]=0
# Mixed Array data[2][3][3][0]=1
# Mixed Array data[2][3][2][2]=0
# Mixed Array data[2][3][2][1]=1
# Mixed Array data[2][3][2][0]=0
# Mixed Array data[2][3][1][2]=1
# Mixed Array data[2][3][1][1]=1
# Mixed Array data[2][3][1][0]=0
# Mixed Array data[2][3][0][2]=1
# Mixed Array data[2][3][0][1]=0
# Mixed Array data[2][3][0][0]=0
# Mixed Array data[2][2][3][2]=0
# Mixed Array data[2][2][3][1]=1
# Mixed Array data[2][2][3][0]=0
# Mixed Array data[2][2][2][2]=1
# Mixed Array data[2][2][2][1]=1
# Mixed Array data[2][2][2][0]=1
# Mixed Array data[2][2][1][2]=1
# Mixed Array data[2][2][1][1]=0
# Mixed Array data[2][2][1][0]=0
# Mixed Array data[2][2][0][2]=0
# Mixed Array data[2][2][0][1]=0
# Mixed Array data[2][2][0][0]=1
# Mixed Array data[2][1][3][2]=0
# Mixed Array data[2][1][3][1]=1
# Mixed Array data[2][1][3][0]=1
# Mixed Array data[2][1][2][2]=1
# Mixed Array data[2][1][2][1]=1
# Mixed Array data[2][1][2][0]=1
# Mixed Array data[2][1][1][2]=0
# Mixed Array data[2][1][1][1]=0
# Mixed Array data[2][1][1][0]=1
# Mixed Array data[2][1][0][2]=1
# Mixed Array data[2][1][0][1]=1
# Mixed Array data[2][1][0][0]=0
# Mixed Array data[2][0][3][2]=0
# Mixed Array data[2][0][3][1]=0
# Mixed Array data[2][0][3][0]=0
# Mixed Array data[2][0][2][2]=0
# Mixed Array data[2][0][2][1]=1
# Mixed Array data[2][0][2][0]=0
# Mixed Array data[2][0][1][2]=0
# Mixed Array data[2][0][1][1]=1
# Mixed Array data[2][0][1][0]=1
# Mixed Array data[2][0][0][2]=0
# Mixed Array data[2][0][0][1]=0
# Mixed Array data[2][0][0][0]=0
# Mixed Array data[1][4][3][2]=0
# Mixed Array data[1][4][3][1]=0
# Mixed Array data[1][4][3][0]=1
# Mixed Array data[1][4][2][2]=1
# Mixed Array data[1][4][2][1]=1
# Mixed Array data[1][4][2][0]=1
# Mixed Array data[1][4][1][2]=1
# Mixed Array data[1][4][1][1]=0
# Mixed Array data[1][4][1][0]=0
# Mixed Array data[1][4][0][2]=1
# Mixed Array data[1][4][0][1]=1
# Mixed Array data[1][4][0][0]=1
# Mixed Array data[1][3][3][2]=0
# Mixed Array data[1][3][3][1]=0
# Mixed Array data[1][3][3][0]=1
# Mixed Array data[1][3][2][2]=1
# Mixed Array data[1][3][2][1]=0
# Mixed Array data[1][3][2][0]=1
# Mixed Array data[1][3][1][2]=1
# Mixed Array data[1][3][1][1]=0
# Mixed Array data[1][3][1][0]=1
# Mixed Array data[1][3][0][2]=1
# Mixed Array data[1][3][0][1]=1
# Mixed Array data[1][3][0][0]=0
# Mixed Array data[1][2][3][2]=1
# Mixed Array data[1][2][3][1]=1
# Mixed Array data[1][2][3][0]=0
# Mixed Array data[1][2][2][2]=0
# Mixed Array data[1][2][2][1]=0
# Mixed Array data[1][2][2][0]=0
# Mixed Array data[1][2][1][2]=1
# Mixed Array data[1][2][1][1]=1
# Mixed Array data[1][2][1][0]=0
# Mixed Array data[1][2][0][2]=0
# Mixed Array data[1][2][0][1]=1
# Mixed Array data[1][2][0][0]=1
# Mixed Array data[1][1][3][2]=1
# Mixed Array data[1][1][3][1]=1
# Mixed Array data[1][1][3][0]=1
# Mixed Array data[1][1][2][2]=0
# Mixed Array data[1][1][2][1]=1
# Mixed Array data[1][1][2][0]=1
# Mixed Array data[1][1][1][2]=1
# Mixed Array data[1][1][1][1]=0
# Mixed Array data[1][1][1][0]=0
# Mixed Array data[1][1][0][2]=0
# Mixed Array data[1][1][0][1]=0
# Mixed Array data[1][1][0][0]=0
# Mixed Array data[1][0][3][2]=0
# Mixed Array data[1][0][3][1]=0
# Mixed Array data[1][0][3][0]=1
# Mixed Array data[1][0][2][2]=1
# Mixed Array data[1][0][2][1]=1
# Mixed Array data[1][0][2][0]=1
# Mixed Array data[1][0][1][2]=1
# Mixed Array data[1][0][1][1]=0
# Mixed Array data[1][0][1][0]=1
# Mixed Array data[1][0][0][2]=1
# Mixed Array data[1][0][0][1]=0
# Mixed Array data[1][0][0][0]=0
# Mixed Array data[0][4][3][2]=1
# Mixed Array data[0][4][3][1]=1
# Mixed Array data[0][4][3][0]=0
# Mixed Array data[0][4][2][2]=1
# Mixed Array data[0][4][2][1]=1
# Mixed Array data[0][4][2][0]=1
# Mixed Array data[0][4][1][2]=1
# Mixed Array data[0][4][1][1]=0
# Mixed Array data[0][4][1][0]=0
# Mixed Array data[0][4][0][2]=0
# Mixed Array data[0][4][0][1]=1
# Mixed Array data[0][4][0][0]=0
# Mixed Array data[0][3][3][2]=0
# Mixed Array data[0][3][3][1]=0
# Mixed Array data[0][3][3][0]=1
# Mixed Array data[0][3][2][2]=1
# Mixed Array data[0][3][2][1]=0
# Mixed Array data[0][3][2][0]=0
# Mixed Array data[0][3][1][2]=1
# Mixed Array data[0][3][1][1]=0
# Mixed Array data[0][3][1][0]=0
# Mixed Array data[0][3][0][2]=0
# Mixed Array data[0][3][0][1]=1
# Mixed Array data[0][3][0][0]=0
# Mixed Array data[0][2][3][2]=0
# Mixed Array data[0][2][3][1]=1
# Mixed Array data[0][2][3][0]=0
# Mixed Array data[0][2][2][2]=1
# Mixed Array data[0][2][2][1]=1
# Mixed Array data[0][2][2][0]=1
# Mixed Array data[0][2][1][2]=1
# Mixed Array data[0][2][1][1]=1
# Mixed Array data[0][2][1][0]=0
# Mixed Array data[0][2][0][2]=0
# Mixed Array data[0][2][0][1]=0
# Mixed Array data[0][2][0][0]=1
# Mixed Array data[0][1][3][2]=0
# Mixed Array data[0][1][3][1]=0
# Mixed Array data[0][1][3][0]=1
# Mixed Array data[0][1][2][2]=1
# Mixed Array data[0][1][2][1]=0
# Mixed Array data[0][1][2][0]=0
# Mixed Array data[0][1][1][2]=0
# Mixed Array data[0][1][1][1]=1
# Mixed Array data[0][1][1][0]=1
# Mixed Array data[0][1][0][2]=0
# Mixed Array data[0][1][0][1]=0
# Mixed Array data[0][1][0][0]=0
# Mixed Array data[0][0][3][2]=1
# Mixed Array data[0][0][3][1]=1
# Mixed Array data[0][0][3][0]=0
# Mixed Array data[0][0][2][2]=0
# Mixed Array data[0][0][2][1]=0
# Mixed Array data[0][0][2][0]=1
# Mixed Array data[0][0][1][2]=0
# Mixed Array data[0][0][1][1]=0
# Mixed Array data[0][0][1][0]=1
# Mixed Array data[0][0][0][2]=0
# Mixed Array data[0][0][0][1]=0
# Mixed Array data[0][0][0][0]=0
