// Code your design here
module repeat_ex;
  initial begin
    repeat(5)begin
      $display("REPEAT LOOP");
    end
  end
endmodule

# REPEAT LOOP
# REPEAT LOOP
# REPEAT LOOP
# REPEAT LOOP
# REPEAT LOOP
